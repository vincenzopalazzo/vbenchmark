module main

import internal

/// Init the benchamarks
fn init_benchamars() {
	internal.init_benchamars()
}

fn main() {
	init_benchamars()
	println('Hello World!')
}
